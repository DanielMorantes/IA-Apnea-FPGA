LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-------------------------------------
ENTITY control_conv IS
	PORT( 	clk						:		IN		STD_LOGIC;
				rst						:		IN		STD_LOGIC;
				
				n_Control_Conv			:		IN		STD_LOGIC; --Enable Control 
				
				Flag_count_RAM			:		IN		STD_LOGIC; --OUT  comparador con 23
				Flag_count_Relu		:		IN		STD_LOGIC; --Flags contadores
				Flag_count_Filtro		:		IN		STD_LOGIC;
				--Flag_countROM_Filtro	:		IN		STD_LOGIC;
				Flag_count_Fin			:		IN		STD_LOGIC;
				
				ena_RAM_1				:		OUT	STD_LOGIC; --Enables RAM's entrada
				ena_RAM_2				:		OUT	STD_LOGIC;
				ena_RAM_3				:		OUT	STD_LOGIC;
				ena_RAM_4				:		OUT	STD_LOGIC;
				ena_RAM_5				:		OUT	STD_LOGIC;
				ena_RAM_6				:		OUT	STD_LOGIC;
				ena_RAM_7				:		OUT	STD_LOGIC;
				ena_RAM_8				:		OUT	STD_LOGIC;
				
				rden						:		OUT	STD_LOGIC; --Enable ROM
					
				enab_reg_ROM_1			:		OUT	STD_LOGIC; --Enables registros ROM
				enab_reg_ROM_2			:		OUT	STD_LOGIC;	
				enab_reg_ROM_3			:		OUT	STD_LOGIC;
				enab_reg_ROM_4			:		OUT	STD_LOGIC;
				enab_reg_ROM_5			:		OUT	STD_LOGIC;
				enab_reg_ROM_6			:		OUT	STD_LOGIC;	
				enab_reg_ROM_7			:		OUT	STD_LOGIC;
				enab_reg_ROM_8			:		OUT	STD_LOGIC;

				reg_raro_rst1			:		OUT	STD_LOGIC; --Resets Registros ROM
				reg_raro_rst2			:		OUT	STD_LOGIC;
				reg_raro_rst3			:		OUT	STD_LOGIC;
				reg_raro_rst4			:		OUT	STD_LOGIC;
				reg_raro_rst5			:		OUT	STD_LOGIC;
				reg_raro_rst6			:		OUT	STD_LOGIC;
				reg_raro_rst7			:		OUT	STD_LOGIC;
				reg_raro_rst8			:		OUT	STD_LOGIC;

				reg_in_ena_1			:		OUT	STD_LOGIC; --Enables registros entrada
				reg_in_ena_2			:		OUT	STD_LOGIC;
				reg_in_ena_3			:		OUT	STD_LOGIC;
				reg_in_ena_4			:		OUT	STD_LOGIC;
				reg_in_ena_5			:		OUT	STD_LOGIC;
				reg_in_ena_6			:		OUT	STD_LOGIC;
				reg_in_ena_7			:		OUT	STD_LOGIC;
				reg_in_ena_8			:		OUT	STD_LOGIC;
		
				reg_in_rst_1			:		OUT	STD_LOGIC; --Resets registros entrada
				reg_in_rst_2			:		OUT	STD_LOGIC;
				reg_in_rst_3			:		OUT	STD_LOGIC;
				reg_in_rst_4			:		OUT	STD_LOGIC;
				reg_in_rst_5			:		OUT	STD_LOGIC;
				reg_in_rst_6			:		OUT	STD_LOGIC;
				reg_in_rst_7			:		OUT	STD_LOGIC;
				reg_in_rst_8			:		OUT	STD_LOGIC;

				reLU_ena					:		OUT	STD_LOGIC; --RELU
				reLU_rst					:		OUT	STD_LOGIC;
		
				reg_Filt_ena			:		OUT	STD_LOGIC; --Registro realimentado
				reg_Filt_rst			:		OUT	STD_LOGIC;

				ctr_count_RAM			:		OUT	STD_LOGIC; --Enables contadores
				ctr_count_Relu			:		OUT	STD_LOGIC;
				ctr_count_Filtro		:		OUT	STD_LOGIC;
				ctr_countROM_Filtro	:		OUT	STD_LOGIC;
				ctr_count_Fin			:		OUT	STD_LOGIC;
				
				Load_count				:		OUT	STD_LOGIC;
		
				rst_count_RAM			:		OUT	STD_LOGIC; --Resets contadores
				rst_count_Relu			:		OUT	STD_LOGIC;
				rst_count_Filtro		:		OUT	STD_LOGIC;
				rst_countROM_Filtro	:		OUT	STD_LOGIC;
				rst_count_Fin			:		OUT	STD_LOGIC;
				n_Max_Pooling			:		OUT	STD_LOGIC;
				n_8byt					:		OUT	STD_LOGIC
				
				);												
END ENTITY;
--------------------------------------
ARCHITECTURE behavioral OF control_conv	IS

	TYPE estados IS (CERO,UNO,UNOYMEDIO,UNOTRESCUARTOS,DOS,ESPERA1,TRES,CUATRO,CUATROYMEDIO,CUATROTRESCUARTOS,CINCO,ESPERA2,SEIS,SIETE,SIETEYMEDIO,SIETETRESCUARTOS,OCHO,ESPERA3,NUEVE,DIEZ,DIEZYMEDIO,DIEZTRESCUARTOS,ONCE,ESPERA4,DOCE,TRECE,CATORCE,QUINCE,DIECISEIS,DIECISIETE);
	SIGNAL state: estados; 
	
BEGIN


	PROCESS (rst,clk,n_Control_Conv)
	BEGIN
			IF(rst='1') THEN
					state <= CERO;
			ELSIF(rising_edge(clk)) THEN
				IF ((rst= '0')) THEN
						CASE state IS
								WHEN	CERO =>
											ena_RAM_1				 <= '0'; --Enables entrada
											ena_RAM_2				 <= '0';
											ena_RAM_3				 <= '0';
											ena_RAM_4				 <= '0';
											ena_RAM_5				 <= '0';
											ena_RAM_6				 <= '0';
											ena_RAM_7				 <= '0';
											ena_RAM_8				 <= '0';
											rden						 <= '0'; --Enables ROMS
											enab_reg_ROM_1			 <= '0'; --Enables registros ROM
											enab_reg_ROM_2			 <= '0';	
											enab_reg_ROM_3			 <= '0';
											enab_reg_ROM_4			 <= '0';
											enab_reg_ROM_5			 <= '0';
											enab_reg_ROM_6			 <= '0';	
											enab_reg_ROM_7			 <= '0';
											enab_reg_ROM_8			 <= '0';
											reg_raro_rst1			 <= '0'; --Resets Registros ROM
											reg_raro_rst2			 <= '0';
											reg_raro_rst3			 <= '0';
											reg_raro_rst4			 <= '0';
											reg_raro_rst5			 <= '0';
											reg_raro_rst6			 <= '0';
											reg_raro_rst7			 <= '0';
											reg_raro_rst8			 <= '0';
											reg_in_ena_1			 <= '0'; --Enables registros entrada
											reg_in_ena_2			 <= '0';
											reg_in_ena_3			 <= '0';
											reg_in_ena_4			 <= '0';
											reg_in_ena_5			 <= '0';
											reg_in_ena_6			 <= '0';
											reg_in_ena_7			 <= '0';
											reg_in_ena_8			 <= '0';
											reg_in_rst_1			 <= '0'; --Resets registros entrada
											reg_in_rst_2			 <= '0';
											reg_in_rst_3			 <= '0';
											reg_in_rst_4			 <= '0';
											reg_in_rst_5			 <= '0';
											reg_in_rst_6			 <= '0';
											reg_in_rst_7			 <= '0';
											reg_in_rst_8			 <= '0';
											reLU_ena					 <= '0'; --RELU
											reLU_rst					 <= '0';
											reg_Filt_ena			 <= '0'; --Registro realimentado
											reg_Filt_rst			 <= '0';
											ctr_count_RAM			 <= '0'; --Enables contadores
											ctr_count_Relu			 <= '0';
											ctr_count_Filtro		 <= '0';
											ctr_countROM_Filtro	 <= '0';
											ctr_count_Fin			 <= '0';
											Load_count			    <= '0';
											rst_count_RAM			 <= '0'; --Resets contadores
											rst_count_Relu			 <= '0';
											rst_count_Filtro		 <= '0';
											rst_countROM_Filtro	 <= '0';
											rst_count_Fin			 <= '0';
											n_Max_Pooling			 <= '0';
											n_8byt					 <= '0';
										IF (n_Control_Conv = '1') THEN			
												state <= UNO;
										 ELSE
												state <= CERO;
										 END IF;
																			    										 
							   WHEN	UNO =>
											ena_RAM_1				 <= '1'; --Enables entrada
											ena_RAM_2				 <= '1';
											ena_RAM_3				 <= '1';
											ena_RAM_4				 <= '1';
											ena_RAM_5				 <= '1';
											ena_RAM_6				 <= '0';
											ena_RAM_7				 <= '0';
											ena_RAM_8				 <= '0';
											rden						 <= '1'; --Enables ROMS (SERIA SOLO UNO XD)
											enab_reg_ROM_1			 <= '0'; --Enables registros ROM
											enab_reg_ROM_2			 <= '0';	
											enab_reg_ROM_3			 <= '0';
											enab_reg_ROM_4			 <= '0';
											enab_reg_ROM_5			 <= '0';
											enab_reg_ROM_6			 <= '0';	
											enab_reg_ROM_7			 <= '0';
											enab_reg_ROM_8			 <= '0';
											reg_raro_rst1			 <= '0'; --Resets Registros ROM
											reg_raro_rst2			 <= '0';
											reg_raro_rst3			 <= '0';
											reg_raro_rst4			 <= '0';
											reg_raro_rst5			 <= '0';
											reg_raro_rst6			 <= '1';
											reg_raro_rst7			 <= '1';
											reg_raro_rst8			 <= '1';
											reg_in_ena_1			 <= '0'; --Enables registros entrada
											reg_in_ena_2			 <= '0';
											reg_in_ena_3			 <= '0';
											reg_in_ena_4			 <= '0';
											reg_in_ena_5			 <= '0';
											reg_in_ena_6			 <= '0';
											reg_in_ena_7			 <= '0';
											reg_in_ena_8			 <= '0';
											reg_in_rst_1			 <= '0'; --Resets registros entrada
											reg_in_rst_2			 <= '0';
											reg_in_rst_3			 <= '0';
											reg_in_rst_4			 <= '0';
											reg_in_rst_5			 <= '0';
											reg_in_rst_6			 <= '1';
											reg_in_rst_7			 <= '1';
											reg_in_rst_8			 <= '1';
											reLU_ena					 <= '0'; --RELU
											reLU_rst					 <= '0';
											reg_Filt_ena			 <= '0'; --Registro realimentado
											reg_Filt_rst			 <= '0';
											ctr_count_RAM			 <= '0'; --Enables contadores
											ctr_count_Relu			 <= '1';
											ctr_count_Filtro		 <= '0';
											ctr_countROM_Filtro	 <= '0';
											ctr_count_Fin			 <= '0';
											Load_count			    <= '0';
											rst_count_RAM			 <= '0'; --Resets contadores
											rst_count_Relu			 <= '0';
											rst_count_Filtro		 <= '0';
											rst_countROM_Filtro	 <= '0';
											rst_count_Fin			 <= '0';
											n_Max_Pooling			 <= '0';	
											n_8byt					 <= '0';					
										 state <= UNOYMEDIO;
										 
								WHEN  UNOYMEDIO =>
											ena_RAM_1				 <= '0'; --Enables entrada
											ena_RAM_2				 <= '0';
											ena_RAM_3				 <= '0';
											ena_RAM_4				 <= '0';
											ena_RAM_5				 <= '0';
											ena_RAM_6				 <= '0';
											ena_RAM_7				 <= '0';
											ena_RAM_8				 <= '0';
											rden						 <= '0'; --Enable ROM
											enab_reg_ROM_1			 <= '1'; --Enables registros ROM
											enab_reg_ROM_2			 <= '1';	
											enab_reg_ROM_3			 <= '1';
											enab_reg_ROM_4			 <= '1';
											enab_reg_ROM_5			 <= '1';
											enab_reg_ROM_6			 <= '0';	
											enab_reg_ROM_7			 <= '0';
											enab_reg_ROM_8			 <= '0';
											reg_raro_rst1			 <= '0'; --Resets Registros ROM
											reg_raro_rst2			 <= '0';
											reg_raro_rst3			 <= '0';
											reg_raro_rst4			 <= '0';
											reg_raro_rst5			 <= '0';
											reg_raro_rst6			 <= '0';
											reg_raro_rst7			 <= '0';
											reg_raro_rst8			 <= '0';
											reg_in_ena_1			 <= '1'; --Enables registros entrada
											reg_in_ena_2			 <= '1';
											reg_in_ena_3			 <= '1';
											reg_in_ena_4			 <= '1';
											reg_in_ena_5			 <= '1';
											reg_in_ena_6			 <= '0';
											reg_in_ena_7			 <= '0';
											reg_in_ena_8			 <= '0';
											reg_in_rst_1			 <= '0'; --Resets registros entrada
											reg_in_rst_2			 <= '0';
											reg_in_rst_3			 <= '0';
											reg_in_rst_4			 <= '0';
											reg_in_rst_5			 <= '0';
											reg_in_rst_6			 <= '0';
											reg_in_rst_7			 <= '0';
											reg_in_rst_8			 <= '0';
											reLU_ena					 <= '0'; --RELU
											reLU_rst					 <= '0';
											reg_Filt_ena			 <= '0'; --Registro realimentado
											reg_Filt_rst			 <= '0';
											ctr_count_RAM			 <= '0'; --Enables contadores
											ctr_count_Relu			 <= '0';
											ctr_count_Filtro		 <= '0';
											ctr_countROM_Filtro	 <= '0';
											ctr_count_Fin			 <= '0';
											Load_count			    <= '0';
											rst_count_RAM			 <= '0'; --Resets contadores
											rst_count_Relu			 <= '0';
											rst_count_Filtro		 <= '0';
											rst_countROM_Filtro	 <= '0';
											rst_count_Fin			 <= '0';	
											n_Max_Pooling			 <= '0';
											n_8byt					 <= '0';
										 state <= UNOTRESCUARTOS;
								
								WHEN	UNOTRESCUARTOS =>
											ena_RAM_1				 <= '0'; --Enables entrada
											ena_RAM_2				 <= '0';
											ena_RAM_3				 <= '0';
											ena_RAM_4				 <= '0';
											ena_RAM_5				 <= '0';
											ena_RAM_6				 <= '0';
											ena_RAM_7				 <= '0';
											ena_RAM_8				 <= '0';
											rden						 <= '0'; --Enables ROMS (SERIA SOLO UNO XD)
											enab_reg_ROM_1			 <= '0'; --Enables registros ROM
											enab_reg_ROM_2			 <= '0';	
											enab_reg_ROM_3			 <= '0';
											enab_reg_ROM_4			 <= '0';
											enab_reg_ROM_5			 <= '0';
											enab_reg_ROM_6			 <= '0';
											enab_reg_ROM_7			 <= '0';
											enab_reg_ROM_8			 <= '0';
											reg_raro_rst1			 <= '0'; --Resets Registros ROM
											reg_raro_rst2			 <= '0';
											reg_raro_rst3			 <= '0';
											reg_raro_rst4			 <= '0';
											reg_raro_rst5			 <= '0';
											reg_raro_rst6			 <= '0';
											reg_raro_rst7			 <= '0';
											reg_raro_rst8			 <= '0';
											reg_in_ena_1			 <= '0'; --Enables registros entrada
											reg_in_ena_2			 <= '0';
											reg_in_ena_3			 <= '0';
											reg_in_ena_4			 <= '0';
											reg_in_ena_5			 <= '0';
											reg_in_ena_6			 <= '0';
											reg_in_ena_7			 <= '0';
											reg_in_ena_8			 <= '0';
											reg_in_rst_1			 <= '0'; --Resets registros entrada
											reg_in_rst_2			 <= '0';
											reg_in_rst_3			 <= '0';
											reg_in_rst_4			 <= '0';
											reg_in_rst_5			 <= '0';
											reg_in_rst_6			 <= '0';
											reg_in_rst_7			 <= '0';
											reg_in_rst_8			 <= '0';
											reLU_ena					 <= '0'; --RELU
											reLU_rst					 <= '0';
											reg_Filt_ena			 <= '1'; --Registro realimentado
											reg_Filt_rst			 <= '0';
											ctr_count_RAM			 <= '0'; --Enables contadores
											ctr_count_Relu			 <= '0';
											ctr_count_Filtro		 <= '0';
											ctr_countROM_Filtro	 <= '0';
											ctr_count_Fin			 <= '0';
											Load_count			    <= '0';
											rst_count_RAM			 <= '0'; --Resets contadores
											rst_count_Relu			 <= '0';
											rst_count_Filtro		 <= '0';
											rst_countROM_Filtro	 <= '0';
											rst_count_Fin			 <= '0';
											n_Max_Pooling			 <= '0';	
											n_8byt					 <= '0';					
										 state <= DOS;
					
								WHEN	DOS =>
											ena_RAM_1				 <= '0'; --Enables entrada
											ena_RAM_2				 <= '0';
											ena_RAM_3				 <= '0';
											ena_RAM_4				 <= '0';
											ena_RAM_5				 <= '0';
											ena_RAM_6				 <= '0';
											ena_RAM_7				 <= '0';
											ena_RAM_8				 <= '0';
											rden						 <= '0'; --Enables ROM
											enab_reg_ROM_1			 <= '0'; --Enables registros ROM
											enab_reg_ROM_2			 <= '0';	
											enab_reg_ROM_3			 <= '0';
											enab_reg_ROM_4			 <= '0';
											enab_reg_ROM_5			 <= '0';
											enab_reg_ROM_6			 <= '0';	
											enab_reg_ROM_7			 <= '0';
											enab_reg_ROM_8			 <= '0';
											reg_raro_rst1			 <= '0'; --Resets Registros ROM
											reg_raro_rst2			 <= '0';
											reg_raro_rst3			 <= '0';
											reg_raro_rst4			 <= '0';
											reg_raro_rst5			 <= '0';
											reg_raro_rst6			 <= '0';
											reg_raro_rst7			 <= '0';
											reg_raro_rst8			 <= '0';
											reg_in_ena_1			 <= '0'; --Enables registros entrada
											reg_in_ena_2			 <= '0';
											reg_in_ena_3			 <= '0';
											reg_in_ena_4			 <= '0';
											reg_in_ena_5			 <= '0';
											reg_in_ena_6			 <= '0';
											reg_in_ena_7			 <= '0';
											reg_in_ena_8			 <= '0';
											reg_in_rst_1			 <= '0'; --Resets registros entrada
											reg_in_rst_2			 <= '0';
											reg_in_rst_3			 <= '0';
											reg_in_rst_4			 <= '0';
											reg_in_rst_5			 <= '0';
											reg_in_rst_6			 <= '0';
											reg_in_rst_7			 <= '0';
											reg_in_rst_8			 <= '0';
											reLU_ena					 <= '0'; --RELU
											reLU_rst					 <= '0';
											reg_Filt_ena			 <= '0'; --Registro realimentado
											reg_Filt_rst			 <= '0';
											ctr_count_RAM			 <= '0'; --Enables contadores
											ctr_count_Relu			 <= '0';
											ctr_count_Filtro		 <= '0';
											ctr_countROM_Filtro	 <= '0';
											ctr_count_Fin			 <= '0';
											Load_count			    <= '0';
											rst_count_RAM			 <= '0'; --Resets contadores
											rst_count_Relu			 <= '0';
											rst_count_Filtro		 <= '0';
											rst_countROM_Filtro	 <= '0';
											rst_count_Fin			 <= '0';
											n_Max_Pooling			 <= '1';
											n_8byt					 <= '0';	
										 IF (Flag_count_Relu = '1') THEN			
												state <= ESPERA1;
										 ELSIF (Flag_count_Relu = '0') THEN
												state <= UNO;
										 ELSE
												state <= DOS;
										 END IF;
										 
								WHEN	ESPERA1 =>
											ena_RAM_1				 <= '0'; --Enables entrada
											ena_RAM_2				 <= '0';
											ena_RAM_3				 <= '0';
											ena_RAM_4				 <= '0';
											ena_RAM_5				 <= '0';
											ena_RAM_6				 <= '0';
											ena_RAM_7				 <= '0';
											ena_RAM_8				 <= '0';
											rden						 <= '0'; --Enables ROMS (SERIA SOLO UNO XD)
											enab_reg_ROM_1			 <= '0'; --Enables registros ROM
											enab_reg_ROM_2			 <= '0';	
											enab_reg_ROM_3			 <= '0';
											enab_reg_ROM_4			 <= '0';
											enab_reg_ROM_5			 <= '0';
											enab_reg_ROM_6			 <= '0';	
											enab_reg_ROM_7			 <= '0';
											enab_reg_ROM_8			 <= '0';
											reg_raro_rst1			 <= '0'; --Resets Registros ROM
											reg_raro_rst2			 <= '0';
											reg_raro_rst3			 <= '0';
											reg_raro_rst4			 <= '0';
											reg_raro_rst5			 <= '0';
											reg_raro_rst6			 <= '0';
											reg_raro_rst7			 <= '0';
											reg_raro_rst8			 <= '0';
											reg_in_ena_1			 <= '0'; --Enables registros entrada
											reg_in_ena_2			 <= '0';
											reg_in_ena_3			 <= '0';
											reg_in_ena_4			 <= '0';
											reg_in_ena_5			 <= '0';
											reg_in_ena_6			 <= '0';
											reg_in_ena_7			 <= '0';
											reg_in_ena_8			 <= '0';
											reg_in_rst_1			 <= '0'; --Resets registros entrada
											reg_in_rst_2			 <= '0';
											reg_in_rst_3			 <= '0';
											reg_in_rst_4			 <= '0';
											reg_in_rst_5			 <= '0';
											reg_in_rst_6			 <= '0';
											reg_in_rst_7			 <= '0';
											reg_in_rst_8			 <= '0';
											reLU_ena					 <= '1'; --RELU
											reLU_rst					 <= '0';
											reg_Filt_ena			 <= '0'; --Registro realimentado
											reg_Filt_rst			 <= '0';
											ctr_count_RAM			 <= '0'; --Enables contadores
											ctr_count_Relu			 <= '1';
											ctr_count_Filtro		 <= '0';
											ctr_countROM_Filtro	 <= '0';
											ctr_count_Fin			 <= '0';
											Load_count			    <= '0';
											rst_count_RAM			 <= '0'; --Resets contadores
											rst_count_Relu			 <= '1';
											rst_count_Filtro		 <= '0';
											rst_countROM_Filtro	 <= '0';
											rst_count_Fin			 <= '0';
											n_Max_Pooling			 <= '0';	
											n_8byt					 <= '0';					
										 state <= TRES;
								
								WHEN  TRES =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enables ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '1';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';
									n_8byt					 <= '1';	
									state <= CUATRO;
										
								WHEN	CUATRO =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '1';
									ena_RAM_3				 <= '1';
									ena_RAM_4				 <= '1';
									ena_RAM_5				 <= '1';
									ena_RAM_6				 <= '1';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '1'; --Enables ROMS (SERIA SOLO UNO XD)
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '1'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '1';
									reg_raro_rst8			 <= '1';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '1'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '1';
									reg_in_rst_8			 <= '1';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '1';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';	
									n_Max_Pooling			 <= '0';
									n_8byt					 <= '0';	
									state <= CUATROYMEDIO;
										 
								WHEN  CUATROYMEDIO =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enable ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '1';	
									enab_reg_ROM_3			 <= '1';
									enab_reg_ROM_4			 <= '1';
									enab_reg_ROM_5			 <= '1';
									enab_reg_ROM_6			 <= '1';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '1';
									reg_in_ena_3			 <= '1';
									reg_in_ena_4			 <= '1';
									reg_in_ena_5			 <= '1';
									reg_in_ena_6			 <= '1';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';
									n_8byt					 <= '0';	
									state <= CUATROTRESCUARTOS;
								
								WHEN  CUATROTRESCUARTOS =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enable ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '1'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';
									n_8byt					 <= '0';	
									state <= CINCO;
						
								WHEN	CINCO =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enables ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0'; 
										 IF (Flag_count_Relu = '1') THEN	
													state <= ESPERA2;
										 ELSIF (Flag_count_Relu = '0') THEN
												state <= CUATRO;
										 ELSE
												state <= CINCO;
										 END IF;
										 
								WHEN	ESPERA2 =>
											ena_RAM_1				 <= '0'; --Enables entrada
											ena_RAM_2				 <= '0';
											ena_RAM_3				 <= '0';
											ena_RAM_4				 <= '0';
											ena_RAM_5				 <= '0';
											ena_RAM_6				 <= '0';
											ena_RAM_7				 <= '0';
											ena_RAM_8				 <= '0';
											rden						 <= '0'; --Enables ROMS (SERIA SOLO UNO XD)
											enab_reg_ROM_1			 <= '0'; --Enables registros ROM
											enab_reg_ROM_2			 <= '0';	
											enab_reg_ROM_3			 <= '0';
											enab_reg_ROM_4			 <= '0';
											enab_reg_ROM_5			 <= '0';
											enab_reg_ROM_6			 <= '0';	
											enab_reg_ROM_7			 <= '0';
											enab_reg_ROM_8			 <= '0';
											reg_raro_rst1			 <= '0'; --Resets Registros ROM
											reg_raro_rst2			 <= '0';
											reg_raro_rst3			 <= '0';
											reg_raro_rst4			 <= '0';
											reg_raro_rst5			 <= '0';
											reg_raro_rst6			 <= '0';
											reg_raro_rst7			 <= '0';
											reg_raro_rst8			 <= '0';
											reg_in_ena_1			 <= '0'; --Enables registros entrada
											reg_in_ena_2			 <= '0';
											reg_in_ena_3			 <= '0';
											reg_in_ena_4			 <= '0';
											reg_in_ena_5			 <= '0';
											reg_in_ena_6			 <= '0';
											reg_in_ena_7			 <= '0';
											reg_in_ena_8			 <= '0';
											reg_in_rst_1			 <= '0'; --Resets registros entrada
											reg_in_rst_2			 <= '0';
											reg_in_rst_3			 <= '0';
											reg_in_rst_4			 <= '0';
											reg_in_rst_5			 <= '0';
											reg_in_rst_6			 <= '0';
											reg_in_rst_7			 <= '0';
											reg_in_rst_8			 <= '0';
											reLU_ena					 <= '1'; --RELU
											reLU_rst					 <= '0';
											reg_Filt_ena			 <= '0'; --Registro realimentado
											reg_Filt_rst			 <= '0';
											ctr_count_RAM			 <= '0'; --Enables contadores
											ctr_count_Relu			 <= '0';
											ctr_count_Filtro		 <= '0';
											ctr_countROM_Filtro	 <= '0';
											ctr_count_Fin			 <= '0';
											Load_count			    <= '0';
											rst_count_RAM			 <= '0'; --Resets contadores
											rst_count_Relu			 <= '1';
											rst_count_Filtro		 <= '0';
											rst_countROM_Filtro	 <= '0';
											rst_count_Fin			 <= '0';
											n_Max_Pooling			 <= '0';	
											n_8byt					 <= '0';					
										 state <= SEIS; 
								
								WHEN  SEIS =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enables ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '1';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';
									n_8byt					 <= '1';	
									state <= SIETE;
										 
								WHEN	SIETE =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '1';
									ena_RAM_4				 <= '1';
									ena_RAM_5				 <= '1';
									ena_RAM_6				 <= '1';
									ena_RAM_7				 <= '1';
									ena_RAM_8				 <= '0';
									rden						 <= '1'; --Enables ROMS (SERIA SOLO UNO XD)
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '1'; --Resets Registros ROM
									reg_raro_rst2			 <= '1';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '1';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '1'; --Resets registros entrada
									reg_in_rst_2			 <= '1';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '1';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '1';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';	
									n_8byt					 <= '0';				
									state <= SIETEYMEDIO;
										 
								WHEN  SIETEYMEDIO =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enable ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '1';
									enab_reg_ROM_4			 <= '1';
									enab_reg_ROM_5			 <= '1';
									enab_reg_ROM_6			 <= '1';	
									enab_reg_ROM_7			 <= '1';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '1';
									reg_in_ena_4			 <= '1';
									reg_in_ena_5			 <= '1';
									reg_in_ena_6			 <= '1';
									reg_in_ena_7			 <= '1';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores FALTA VALOR INICIO Y LOAD
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';
									n_8byt					 <= '0';
									state <= SIETETRESCUARTOS;
										 
								WHEN  SIETETRESCUARTOS =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enable ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '1'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';
									n_8byt					 <= '0';	
									state <= OCHO;
								
								WHEN	OCHO =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enables ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';
										 IF (Flag_count_Relu = '1') THEN		
												state <= ESPERA3;
										 ELSIF (Flag_count_Relu = '0') THEN
												state <= SIETE;
										 ELSE
												state <= OCHO;
										 END IF;
										 
								WHEN	ESPERA3 =>
											ena_RAM_1				 <= '0'; --Enables entrada
											ena_RAM_2				 <= '0';
											ena_RAM_3				 <= '0';
											ena_RAM_4				 <= '0';
											ena_RAM_5				 <= '0';
											ena_RAM_6				 <= '0';
											ena_RAM_7				 <= '0';
											ena_RAM_8				 <= '0';
											rden						 <= '0'; --Enables ROMS (SERIA SOLO UNO XD)
											enab_reg_ROM_1			 <= '0'; --Enables registros ROM
											enab_reg_ROM_2			 <= '0';	
											enab_reg_ROM_3			 <= '0';
											enab_reg_ROM_4			 <= '0';
											enab_reg_ROM_5			 <= '0';
											enab_reg_ROM_6			 <= '0';	
											enab_reg_ROM_7			 <= '0';
											enab_reg_ROM_8			 <= '0';
											reg_raro_rst1			 <= '0'; --Resets Registros ROM
											reg_raro_rst2			 <= '0';
											reg_raro_rst3			 <= '0';
											reg_raro_rst4			 <= '0';
											reg_raro_rst5			 <= '0';
											reg_raro_rst6			 <= '0';
											reg_raro_rst7			 <= '0';
											reg_raro_rst8			 <= '0';
											reg_in_ena_1			 <= '0'; --Enables registros entrada
											reg_in_ena_2			 <= '0';
											reg_in_ena_3			 <= '0';
											reg_in_ena_4			 <= '0';
											reg_in_ena_5			 <= '0';
											reg_in_ena_6			 <= '0';
											reg_in_ena_7			 <= '0';
											reg_in_ena_8			 <= '0';
											reg_in_rst_1			 <= '0'; --Resets registros entrada
											reg_in_rst_2			 <= '0';
											reg_in_rst_3			 <= '0';
											reg_in_rst_4			 <= '0';
											reg_in_rst_5			 <= '0';
											reg_in_rst_6			 <= '0';
											reg_in_rst_7			 <= '0';
											reg_in_rst_8			 <= '0';
											reLU_ena					 <= '1'; --RELU
											reLU_rst					 <= '0';
											reg_Filt_ena			 <= '0'; --Registro realimentado
											reg_Filt_rst			 <= '0';
											ctr_count_RAM			 <= '0'; --Enables contadores
											ctr_count_Relu			 <= '0';
											ctr_count_Filtro		 <= '0';
											ctr_countROM_Filtro	 <= '0';
											ctr_count_Fin			 <= '0';
											Load_count			    <= '0';
											rst_count_RAM			 <= '0'; --Resets contadores
											rst_count_Relu			 <= '1';
											rst_count_Filtro		 <= '0';
											rst_countROM_Filtro	 <= '0';
											rst_count_Fin			 <= '0';
											n_Max_Pooling			 <= '0';	
											n_8byt					 <= '0';					
										 state <= NUEVE; 		
									
								WHEN  NUEVE =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enables ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '1';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '1';
									n_8byt					 <= '0';	
									state <= DIEZ;
											
								WHEN	DIEZ =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '1';
									ena_RAM_5				 <= '1';
									ena_RAM_6				 <= '1';
									ena_RAM_7				 <= '1';
									ena_RAM_8				 <= '1';
									rden						 <= '1'; --Enables ROMS (SERIA SOLO UNO XD)
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '1'; --Resets Registros ROM
									reg_raro_rst2			 <= '1';
									reg_raro_rst3			 <= '1';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '1'; --Resets registros entrada
									reg_in_rst_2			 <= '1';
									reg_in_rst_3			 <= '1';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '1';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';					
									n_8byt					 <= '0';	
									state <= DIEZYMEDIO;
										 
								WHEN  DIEZYMEDIO =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enable ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '1';
									enab_reg_ROM_5			 <= '1';
									enab_reg_ROM_6			 <= '1';	
									enab_reg_ROM_7			 <= '1';
									enab_reg_ROM_8			 <= '1';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '1';
									reg_in_ena_5			 <= '1';
									reg_in_ena_6			 <= '1';
									reg_in_ena_7			 <= '1';
									reg_in_ena_8			 <= '1';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores 
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';	
									n_Max_Pooling			 <= '0';	
									state <= DIEZTRESCUARTOS;
								
								WHEN  DIEZTRESCUARTOS =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enable ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '1'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';
									n_8byt					 <= '0';	
									state <= ONCE;
					
								WHEN	ONCE =>
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enables ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';
									n_8byt					 <= '0';
										 IF (Flag_count_Relu = '1') THEN
												state <= ESPERA4;
										 ELSIF (Flag_count_Relu = '0') THEN	
												state <= DIEZ;
										 ELSE
												state <= ONCE;
										 END IF;
										 
								WHEN	ESPERA4 =>
											ena_RAM_1				 <= '0'; --Enables entrada
											ena_RAM_2				 <= '0';
											ena_RAM_3				 <= '0';
											ena_RAM_4				 <= '0';
											ena_RAM_5				 <= '0';
											ena_RAM_6				 <= '0';
											ena_RAM_7				 <= '0';
											ena_RAM_8				 <= '0';
											rden						 <= '0'; --Enables ROMS (SERIA SOLO UNO XD)
											enab_reg_ROM_1			 <= '0'; --Enables registros ROM
											enab_reg_ROM_2			 <= '0';	
											enab_reg_ROM_3			 <= '0';
											enab_reg_ROM_4			 <= '0';
											enab_reg_ROM_5			 <= '0';
											enab_reg_ROM_6			 <= '0';	
											enab_reg_ROM_7			 <= '0';
											enab_reg_ROM_8			 <= '0';
											reg_raro_rst1			 <= '0'; --Resets Registros ROM
											reg_raro_rst2			 <= '0';
											reg_raro_rst3			 <= '0';
											reg_raro_rst4			 <= '0';
											reg_raro_rst5			 <= '0';
											reg_raro_rst6			 <= '0';
											reg_raro_rst7			 <= '0';
											reg_raro_rst8			 <= '0';
											reg_in_ena_1			 <= '0'; --Enables registros entrada
											reg_in_ena_2			 <= '0';
											reg_in_ena_3			 <= '0';
											reg_in_ena_4			 <= '0';
											reg_in_ena_5			 <= '0';
											reg_in_ena_6			 <= '0';
											reg_in_ena_7			 <= '0';
											reg_in_ena_8			 <= '0';
											reg_in_rst_1			 <= '0'; --Resets registros entrada
											reg_in_rst_2			 <= '0';
											reg_in_rst_3			 <= '0';
											reg_in_rst_4			 <= '0';
											reg_in_rst_5			 <= '0';
											reg_in_rst_6			 <= '0';
											reg_in_rst_7			 <= '0';
											reg_in_rst_8			 <= '0';
											reLU_ena					 <= '1'; --RELU
											reLU_rst					 <= '0';
											reg_Filt_ena			 <= '0'; --Registro realimentado
											reg_Filt_rst			 <= '0';
											ctr_count_RAM			 <= '0'; --Enables contadores
											ctr_count_Relu			 <= '0';
											ctr_count_Filtro		 <= '0';
											ctr_countROM_Filtro	 <= '0';
											ctr_count_Fin			 <= '0';
											Load_count			    <= '0';
											rst_count_RAM			 <= '0'; --Resets contadores
											rst_count_Relu			 <= '1';
											rst_count_Filtro		 <= '0';
											rst_countROM_Filtro	 <= '0';
											rst_count_Fin			 <= '0';
											n_Max_Pooling			 <= '0';	
											n_8byt					 <= '0';					
										  state <= DOCE; 
										 
								WHEN  DOCE => 
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enables ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '1';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';
									n_8byt					 <= '1';	
									state <= TRECE;
										 
								WHEN TRECE => 
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enables ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '1';
									Load_count			    <= '0';-- NO SE USA XD
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';
									n_8byt					 <= '1';	
									state <= CATORCE;
										
								WHEN CATORCE => 
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enables ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			 	 <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0'; 
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';
									n_8byt					 <= '0';
										 IF (Flag_count_Fin = '0') THEN
												state <= UNO;
										 ELSIF (Flag_count_Fin = '1') THEN	
												state <= QUINCE;
										 ELSE
												state <= CATORCE;
										 END IF;
										 
								WHEN QUINCE => 
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enables ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '1';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '1';
									n_Max_Pooling			 <= '0';
									n_8byt					 <= '0';
									state <= DIECISEIS;
									
								WHEN DIECISEIS => 
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enables ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '0'; --Resets Registros ROM
									reg_raro_rst2			 <= '0';
									reg_raro_rst3			 <= '0';
									reg_raro_rst4			 <= '0';
									reg_raro_rst5			 <= '0';
									reg_raro_rst6			 <= '0';
									reg_raro_rst7			 <= '0';
									reg_raro_rst8			 <= '0';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '0'; --Resets registros entrada
									reg_in_rst_2			 <= '0';
									reg_in_rst_3			 <= '0';
									reg_in_rst_4			 <= '0';
									reg_in_rst_5			 <= '0';
									reg_in_rst_6			 <= '0';
									reg_in_rst_7			 <= '0';
									reg_in_rst_8			 <= '0';
									reLU_ena					 <= '0'; --RELU
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			 	 <= '0';
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '0';
									rst_countROM_Filtro	 <= '0'; 
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';
									n_8byt					 <= '0';
										 IF (Flag_count_Filtro = '0') THEN
												state <= UNO;
										 ELSIF (Flag_count_Filtro = '1') THEN	
												state <= DIECISIETE;
										 ELSE
												state <= DIECISEIS;
										 END IF;
								WHEN DIECISIETE => 
									ena_RAM_1				 <= '0'; --Enables entrada
									ena_RAM_2				 <= '0';
									ena_RAM_3				 <= '0';
									ena_RAM_4				 <= '0';
									ena_RAM_5				 <= '0';
									ena_RAM_6				 <= '0';
									ena_RAM_7				 <= '0';
									ena_RAM_8				 <= '0';
									rden						 <= '0'; --Enables ROM
									enab_reg_ROM_1			 <= '0'; --Enables registros ROM
									enab_reg_ROM_2			 <= '0';	
									enab_reg_ROM_3			 <= '0';
									enab_reg_ROM_4			 <= '0';
									enab_reg_ROM_5			 <= '0';
									enab_reg_ROM_6			 <= '0';	
									enab_reg_ROM_7			 <= '0';
									enab_reg_ROM_8			 <= '0';
									reg_raro_rst1			 <= '1'; --Resets Registros ROM
									reg_raro_rst2			 <= '1';
									reg_raro_rst3			 <= '1';
									reg_raro_rst4			 <= '1';
									reg_raro_rst5			 <= '1';
									reg_raro_rst6			 <= '1';
									reg_raro_rst7			 <= '1';
									reg_raro_rst8			 <= '1';
									reg_in_ena_1			 <= '0'; --Enables registros entrada
									reg_in_ena_2			 <= '0';
									reg_in_ena_3			 <= '0';
									reg_in_ena_4			 <= '0';
									reg_in_ena_5			 <= '0';
									reg_in_ena_6			 <= '0';
									reg_in_ena_7			 <= '0';
									reg_in_ena_8			 <= '0';
									reg_in_rst_1			 <= '1'; --Resets registros entrada
									reg_in_rst_2			 <= '1';
									reg_in_rst_3			 <= '1';
									reg_in_rst_4			 <= '1';
									reg_in_rst_5			 <= '1';
									reg_in_rst_6			 <= '1';
									reg_in_rst_7			 <= '1';
									reg_in_rst_8			 <= '1';
									reLU_ena					 <= '0'; --RELU SALIDA SIGUIENTE FILTRO
									reLU_rst					 <= '0';
									reg_Filt_ena			 <= '0'; --Registro realimentado
									reg_Filt_rst			 <= '0';
									ctr_count_RAM			 <= '0'; --Enables contadores
									ctr_count_Relu			 <= '0';
									ctr_count_Filtro		 <= '0';
									ctr_countROM_Filtro	 <= '0';
									ctr_count_Fin			 <= '0';
									Load_count			    <= '0';-- NO SE USA XD
									rst_count_RAM			 <= '0'; --Resets contadores
									rst_count_Relu			 <= '0';
									rst_count_Filtro		 <= '1';
									rst_countROM_Filtro	 <= '0';
									rst_count_Fin			 <= '0';
									n_Max_Pooling			 <= '0';--ACABE TODO
									n_8byt					 <= '0';
									state <= CERO;
									
									
							END CASE;
					END IF;
			END IF;
	END PROCESS;
	
	
END ARCHITECTURE;