-- megafunction wizard: %PARALLEL_ADD%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: parallel_add 

-- ============================================================
-- File Name: Sum1Capa2.vhd
-- Megafunction Name(s):
-- 			parallel_add
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 15.0.0 Build 145 04/22/2015 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus II License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY Sum1Capa2 IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (43 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (43 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (43 DOWNTO 0)
	);
END Sum1Capa2;


ARCHITECTURE SYN OF sum1capa2 IS

--	type ALTERA_MF_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (43 DOWNTO 0);
	SIGNAL sub_wire1	: ALTERA_MF_LOGIC_2D (1 DOWNTO 0, 43 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (43 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (43 DOWNTO 0);

BEGIN
	sub_wire2    <= data0x(43 DOWNTO 0);
	sub_wire0    <= data1x(43 DOWNTO 0);
	sub_wire1(1, 0)    <= sub_wire0(0);
	sub_wire1(1, 1)    <= sub_wire0(1);
	sub_wire1(1, 2)    <= sub_wire0(2);
	sub_wire1(1, 3)    <= sub_wire0(3);
	sub_wire1(1, 4)    <= sub_wire0(4);
	sub_wire1(1, 5)    <= sub_wire0(5);
	sub_wire1(1, 6)    <= sub_wire0(6);
	sub_wire1(1, 7)    <= sub_wire0(7);
	sub_wire1(1, 8)    <= sub_wire0(8);
	sub_wire1(1, 9)    <= sub_wire0(9);
	sub_wire1(1, 10)    <= sub_wire0(10);
	sub_wire1(1, 11)    <= sub_wire0(11);
	sub_wire1(1, 12)    <= sub_wire0(12);
	sub_wire1(1, 13)    <= sub_wire0(13);
	sub_wire1(1, 14)    <= sub_wire0(14);
	sub_wire1(1, 15)    <= sub_wire0(15);
	sub_wire1(1, 16)    <= sub_wire0(16);
	sub_wire1(1, 17)    <= sub_wire0(17);
	sub_wire1(1, 18)    <= sub_wire0(18);
	sub_wire1(1, 19)    <= sub_wire0(19);
	sub_wire1(1, 20)    <= sub_wire0(20);
	sub_wire1(1, 21)    <= sub_wire0(21);
	sub_wire1(1, 22)    <= sub_wire0(22);
	sub_wire1(1, 23)    <= sub_wire0(23);
	sub_wire1(1, 24)    <= sub_wire0(24);
	sub_wire1(1, 25)    <= sub_wire0(25);
	sub_wire1(1, 26)    <= sub_wire0(26);
	sub_wire1(1, 27)    <= sub_wire0(27);
	sub_wire1(1, 28)    <= sub_wire0(28);
	sub_wire1(1, 29)    <= sub_wire0(29);
	sub_wire1(1, 30)    <= sub_wire0(30);
	sub_wire1(1, 31)    <= sub_wire0(31);
	sub_wire1(1, 32)    <= sub_wire0(32);
	sub_wire1(1, 33)    <= sub_wire0(33);
	sub_wire1(1, 34)    <= sub_wire0(34);
	sub_wire1(1, 35)    <= sub_wire0(35);
	sub_wire1(1, 36)    <= sub_wire0(36);
	sub_wire1(1, 37)    <= sub_wire0(37);
	sub_wire1(1, 38)    <= sub_wire0(38);
	sub_wire1(1, 39)    <= sub_wire0(39);
	sub_wire1(1, 40)    <= sub_wire0(40);
	sub_wire1(1, 41)    <= sub_wire0(41);
	sub_wire1(1, 42)    <= sub_wire0(42);
	sub_wire1(1, 43)    <= sub_wire0(43);
	sub_wire1(0, 0)    <= sub_wire2(0);
	sub_wire1(0, 1)    <= sub_wire2(1);
	sub_wire1(0, 2)    <= sub_wire2(2);
	sub_wire1(0, 3)    <= sub_wire2(3);
	sub_wire1(0, 4)    <= sub_wire2(4);
	sub_wire1(0, 5)    <= sub_wire2(5);
	sub_wire1(0, 6)    <= sub_wire2(6);
	sub_wire1(0, 7)    <= sub_wire2(7);
	sub_wire1(0, 8)    <= sub_wire2(8);
	sub_wire1(0, 9)    <= sub_wire2(9);
	sub_wire1(0, 10)    <= sub_wire2(10);
	sub_wire1(0, 11)    <= sub_wire2(11);
	sub_wire1(0, 12)    <= sub_wire2(12);
	sub_wire1(0, 13)    <= sub_wire2(13);
	sub_wire1(0, 14)    <= sub_wire2(14);
	sub_wire1(0, 15)    <= sub_wire2(15);
	sub_wire1(0, 16)    <= sub_wire2(16);
	sub_wire1(0, 17)    <= sub_wire2(17);
	sub_wire1(0, 18)    <= sub_wire2(18);
	sub_wire1(0, 19)    <= sub_wire2(19);
	sub_wire1(0, 20)    <= sub_wire2(20);
	sub_wire1(0, 21)    <= sub_wire2(21);
	sub_wire1(0, 22)    <= sub_wire2(22);
	sub_wire1(0, 23)    <= sub_wire2(23);
	sub_wire1(0, 24)    <= sub_wire2(24);
	sub_wire1(0, 25)    <= sub_wire2(25);
	sub_wire1(0, 26)    <= sub_wire2(26);
	sub_wire1(0, 27)    <= sub_wire2(27);
	sub_wire1(0, 28)    <= sub_wire2(28);
	sub_wire1(0, 29)    <= sub_wire2(29);
	sub_wire1(0, 30)    <= sub_wire2(30);
	sub_wire1(0, 31)    <= sub_wire2(31);
	sub_wire1(0, 32)    <= sub_wire2(32);
	sub_wire1(0, 33)    <= sub_wire2(33);
	sub_wire1(0, 34)    <= sub_wire2(34);
	sub_wire1(0, 35)    <= sub_wire2(35);
	sub_wire1(0, 36)    <= sub_wire2(36);
	sub_wire1(0, 37)    <= sub_wire2(37);
	sub_wire1(0, 38)    <= sub_wire2(38);
	sub_wire1(0, 39)    <= sub_wire2(39);
	sub_wire1(0, 40)    <= sub_wire2(40);
	sub_wire1(0, 41)    <= sub_wire2(41);
	sub_wire1(0, 42)    <= sub_wire2(42);
	sub_wire1(0, 43)    <= sub_wire2(43);
	result    <= sub_wire3(43 DOWNTO 0);

	parallel_add_component : parallel_add
	GENERIC MAP (
		msw_subtract => "NO",
		pipeline => 0,
		representation => "SIGNED",
		result_alignment => "LSB",
		shift => 0,
		size => 2,
		width => 44,
		widthr => 44,
		lpm_type => "parallel_add"
	)
	PORT MAP (
		data => sub_wire1,
		result => sub_wire3
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: MSW_SUBTRACT STRING "NO"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "0"
-- Retrieval info: CONSTANT: REPRESENTATION STRING "SIGNED"
-- Retrieval info: CONSTANT: RESULT_ALIGNMENT STRING "LSB"
-- Retrieval info: CONSTANT: SHIFT NUMERIC "0"
-- Retrieval info: CONSTANT: SIZE NUMERIC "2"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "44"
-- Retrieval info: CONSTANT: WIDTHR NUMERIC "44"
-- Retrieval info: USED_PORT: data0x 0 0 44 0 INPUT NODEFVAL "data0x[43..0]"
-- Retrieval info: USED_PORT: data1x 0 0 44 0 INPUT NODEFVAL "data1x[43..0]"
-- Retrieval info: USED_PORT: result 0 0 44 0 OUTPUT NODEFVAL "result[43..0]"
-- Retrieval info: CONNECT: @data 1 0 44 0 data0x 0 0 44 0
-- Retrieval info: CONNECT: @data 1 1 44 0 data1x 0 0 44 0
-- Retrieval info: CONNECT: result 0 0 44 0 @result 0 0 44 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL Sum1Capa2.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Sum1Capa2.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Sum1Capa2.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Sum1Capa2.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Sum1Capa2_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
