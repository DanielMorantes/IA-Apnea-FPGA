LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-------------------------------------

ENTITY Registro_ROM_6in IS
	PORT( 	clk				:		IN		STD_LOGIC;
				n_Res				:		IN		STD_LOGIC;
				Ena_2				:		IN 	STD_LOGIC;	
				Ena_3				:		IN 	STD_LOGIC;	
				Ena_4				:		IN 	STD_LOGIC;
				Ena_5				:		IN 	STD_LOGIC;
				Ena_6				:		IN 	STD_LOGIC;	
				Registro_IN_3	:		IN		STD_LOGIC_VECTOR (7 DOWNTO 0);
				Registro_IN_4	:		IN		STD_LOGIC_VECTOR (7 DOWNTO 0);
				Registro_IN_5	:		IN		STD_LOGIC_VECTOR (7 DOWNTO 0);
				
				Registro_OUT	:		OUT	STD_LOGIC_VECTOR(7 DOWNTO 0)
	);												
END ENTITY;

-------------------------------------
architecture Registro_Arch of Registro_ROM_6in is
SIGNAL estado: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN

PROCESS (clk, n_Res, Ena_2, Ena_3, Ena_4, Ena_5, Ena_6, Registro_IN_3, Registro_IN_4, Registro_IN_5)
BEGIN 
IF ( n_Res = '1') THEN
	estado <= "00000000";
ELSIF (rising_edge(clk)) THEN
	IF ((Ena_2 = '1') AND (Ena_3 = '1') AND (Ena_4 = '1') AND (Ena_5 = '1') AND (Ena_6 = '1')) THEN
		estado <= Registro_IN_5;	
	ELSIF ((Ena_2 = '0') AND (Ena_3 = '1') AND (Ena_4 = '1') AND (Ena_5 = '1') AND (Ena_6 = '1')) THEN
		estado <= Registro_IN_4;
	ELSIF ((Ena_2 = '0') AND (Ena_3 = '0') AND (Ena_4 = '1') AND (Ena_5 = '1') AND (Ena_6 = '1')) THEN
		estado <= Registro_IN_3;
	ELSE
		estado <= estado;
	END IF;
END IF;

END PROCESS;

Registro_OUT <= estado;


End Registro_Arch;